//-----------------------------------------------------------
//-----------------------------------------------------------
//---------* Next PC Logic Combinational Circuit *-----------
//-----------------------------------------------------------
//-----------------------------------------------------------
//-----------------------------------------------------------
//-----------------------------------------------------------

module NextPCLogic(PCNext, PCPlus4, PC, ImmExt, PCSrc);
       input [63:0] PC, ImmExt;
       input PCSrc;
       output [63:0] PCNext, PCPlus4;
       /* write your code here */
	assign PCPlus4=PC+4;
        assign PCNext=(PCSrc==1)?PC+ ImmExt:PCPlus4;
endmodule
