module add (input [63:0] A1, A2,
output [63:0] Y);
assign Y = A1 + A2;
endmodule

